module nbcac_18di_decoder_core(
		output [17:0] v,
		input [26:1] d
		);

parameter	s1=32'd1,
			s2=32'd150050,
			s3=32'd92736,
			s4=32'd57314,
			s5=32'd35422,
			s6=32'd21892,
			s7=32'd13530,
			s8=32'd8362,
			s9=32'd5168,
			s10=32'd3194,
			s11=32'd1974,
			s12=32'd1220,
			s13=32'd754,
			s14=32'd466,
			s15=32'd288,
			s16=32'd178,
			s17=32'd110,
			s18=32'd68,
			s19=32'd42,
			s20=32'd26,
			s21=32'd16,
			s22=32'd10,
			s23=32'd6,
			s24=32'd4,
			s25=32'd2,
			s26=32'd2;

assign v=s26*d[26]+s25*d[25]+s24*d[24]+s23*d[23]+s22*d[22]+s21*d[21]+s20*d[20]+s19*d[19]+s18*d[18]+s17*d[17]+s16*d[16]+s15*d[15]+s14*d[14]+s13*d[13]+s12*d[12]+s11*d[11]+s10*d[10]+s9*d[9]+s8*d[8]+s7*d[7]+s6*d[6]+s5*d[5]+s4*d[4]+s3*d[3]+s2*d[2]+s1*d[1];

endmodule