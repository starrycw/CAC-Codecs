module IFNS_decoder_10(
    input wire clock,
    input wire rst_n,
    output reg [6:0] dataout,
    input wire [10:1] codein
);

    wire [6:0] dataout_wire;

    decoderIFNS_7di_core core_instance(
        .v(dataout_wire),
        .d10(codein[10]),
        .d9(codein[9]),
        .d8(codein[8]),
        .d7(codein[7]),
        .d6(codein[6]),
        .d5(codein[5]),
        .d4(codein[4]),
        .d3(codein[3]),
        .d2(codein[2]),
        .d1(codein[1])
    );

    //sync
    always @(posedge clock or negedge rst_n) begin
        if (~rst_n) begin
            dataout <= 0;
        end
        else begin
            dataout <= dataout_wire;
        end
    end

endmodule